module ebreak(
    input   [31:0]  inst
);

    always @(*) begin
        if(isnt == )
    end

endmodule